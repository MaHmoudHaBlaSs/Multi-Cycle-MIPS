library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity MDR is
	port (
		clk : in std_logic;
		reg_in   : in std_logic_vector(31 downto 0);
		reg_out  : out std_logic_vector(31 downto 0)
		);
end entity;

architecture reg of MDR is
begin
	process(clk)
	begin
		if(rising_edge(clk)) then
			reg_out <= reg_in;
		end if;
		
	end process;
	
	
end architecture ;